interface intf();
	bit [3:0]a;
	bit [3:0]b;
	bit y1,y2,y3;
endinterface

